module Imem(
    input
        logic [31:0] a,
    output
        logic [31:0] rd
);

// 64KiB memory
logic [31:0] mem[63:0];

initial begin
    mem[1] = 32'b00000000000100000000000010010011; // addi r1, 1(r0)
    mem[2] = 32'b00000000000100000000010000100011; // sb r1, 8(r0)
    mem[3] = 32'b00000000100000000001000100000011; // lh r2, 8(r0)
    mem[4] = 32'b11111111111100000000000000010011; // addi r0, 4095(r0)
    mem[5] = 32'b00000000001000001000000110110011; // add r3, r1, r2
    mem[6] = 32'b11111111000111111111000001101111; // j -16
end

assign rd = mem[a[7:2]];

endmodule

